module Format_Data();


endmodule
